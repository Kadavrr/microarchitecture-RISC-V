module Tract(
	
	);
	
endmodule