module DUT;
endmodule