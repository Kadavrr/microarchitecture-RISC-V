module Tract(
	);
	
endmodule