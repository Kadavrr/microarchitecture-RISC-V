module ImmercialExtension(
	input logic A, 
	output logic ImmExtD);

endmodule